use ieee.std_logic_1164.all;
package date_stamp is
constant revision_date : std_logic_vector(31 downto 0) := X"23042014";
constant revision_time : std_logic_vector(31 downto 0) := X"14382100";
end package date_stamp;
